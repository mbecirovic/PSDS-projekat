library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sonicTest is
    port(clk: in std_logic;
          echo: in std_logic;
          trig: out std_logic;
			 Hex: out std_logic_vector(6 downto 0)
          );
end sonicTest;

architecture s of sonicTest is
	 
	 component sonic is
    port(clk: in std_logic;
          echo: in std_logic;
          trig: out std_logic;
			 adresa_tona: out std_logic_vector(1 downto 0)
          );
	 end component;
		
	component seg27 is
   port(
        i: in unsigned(3 downto 0);
        o : out std_logic_vector(6 downto 0)
    );
	end component;

	signal broj : unsigned(3 downto 0);
	signal adresaT : std_logic_vector(1 downto 0);
	
   begin
	 
	 preuzmiSaSonica : sonic port map(clk,echo,trig,adresaT);
	 ispisNaHex : seg27 port map(broj,Hex);
	 
	 broj <= unsigned("00" & adresaT);
    				
   -- cifra0 <= distanca mod 10;
   -- cifra1 <= distanca /10;
    
    --izlazHex0: FourBit7seg port map(std_logic_vector(to_signed(broj_tipke, 4)), Hex0(0), Hex0(1), Hex0(2), Hex0(3), Hex0(4), Hex0(5), Hex0(6));
   -- izlazHex1: FourBit7seg port map(std_logic_vector(to_signed(cifra0, 4)), Hex1(0), Hex1(1), Hex1(2), Hex1(3), Hex1(4), Hex1(5), Hex1(6));
   -- izlazHex2: FourBit7seg port map(std_logic_vector(to_signed(cifra1, 4)), Hex2(0), Hex2(1), Hex2(2), Hex2(3), Hex2(4), Hex2(5), Hex2(6));

        
end s;